// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7 − 0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs:    LEDR7 − 0 are parallel port outputs from the Nios II system
module DE1_SoC (CLOCK_50, SW, KEY, LEDR, GPIO_0);
	input CLOCK_50;
	input [9:0]  SW;
	input [3:0]  KEY;
	output [9:0]  LEDR;
	inout [35:0] GPIO_0;
	
	reg [25:0] tBase;
	always@(posedge CLOCK_50) tBase <= tBase + 1'b1;
	
	wire receive_reset;
	wire clk = CLOCK_50;
	wire serial_clk;
	wire rst = ~KEY[0];
	wire [7:0] transmitData;
	wire transmitLoad, transmitEnable, charTransmitted, serialDataOut;
	wire [7:0] receiveData;
	wire serialDataIn, charReceived;
	// Following line does not properly synthesize!!!!
	//wire [9:0] transmitInfo = {transmitEnable, transmitLoad, transmitData};
	wire [1:0] status = {charTransmitted, charReceived};
	
	transmit send (.clk(serial_clk), .rst, .load(transmitLoad), .parallelDataIn(transmitData), .transmitEnable, .charSent(charTransmitted), .serialDataOut);
	receive read (.clk(serial_clk), .rst(rst | receive_reset), .serialDataIn, .charReceived, .parallelDataOut(receiveData));

	assign serialDataIn = GPIO_0[0];
	assign GPIO_0[1] = serialDataOut;
	
// Instantiate the Nios II system module generated by the Qsys tool:
	nios_system  NiosII  (
		.clk_clk(clk),
		.serial_clk_clk(serial_clk),
		.reset_reset_n(~rst),
		.switches_export(SW[7:0]),
		.leds_export(LEDR[7:0]),
		.transmit_data_export(transmitData),
		.control_export({receive_reset, transmitEnable, transmitLoad}),
		.receive_data_export(receiveData),
		.status_export(status));

endmodule
